`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    09:11:19 10/03/2012 
// Design Name: 
// Module Name:    seg7 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module seg7(bcd,led,led2);
    input [3:0] bcd;
    output [7:0]led;
	 reg [7:0] led;
	 output [7:0]led2;
	 reg [7:0] led2;
   
	 


always @(bcd)
		
	
			
	
		
		
		case (bcd)       //abcdefg
			0: begin
			led = 8'b00000011;
			led2 = 8'b00000011;
			end
	   	1: begin
			led = 8'b10011111;
			led2 = 8'b00000011;
			end
			2: begin
			led = 8'b00100101;
			led2 = 8'b00000011;
			end
			3: begin
			led = 8'b00001101;
			led2 = 8'b00000011;
			end			
			4: begin
			led = 8'b10011001;
			led2 = 8'b00000011;
			end
			5: led = 8'b01001001;
			5: led2 = 8'b00000011;
			6: led = 8'b01000001;
			6: led2 = 8'b00000011;
			7: led = 8'b00011111;
			7: led2 = 8'b00000011;
			8: led = 8'b00000001;
			8: led2 = 8'b00000011;
			9: led = 8'b00001001;
			9: led2 = 8'b00000011;
	///////////////////////////////////////////		
			
			10: led = 8'b00000011;
	   	10: led2 = 8'b10011111;
			11: led = 8'b10011111;
			11: led2 = 8'b10011111;
			12: led = 8'b00100101;
			12: led2 = 8'b10011111;
			13: led = 8'b00001101;
			13:begin
			led2 = 8'b10011111;
			led = 8'b10011001;
			end
			14: led2 = 8'b10011111;
			15: led = 8'b01001001;
			15: led2 = 8'b10011111;
			16: led = 8'b01000001;
			16: led2 = 8'b10011111;
			17: led = 8'b00011111;
			17: led2 = 8'b10011111;
			18: led = 8'b00000001;
			18: led2 = 8'b10011111;
			19: led = 8'b00001001;
			19: led2 = 8'b10011111;
	//////////////////////////////////////////////////////	
			20: led = 8'b00000011;
	   	20: led2 = 8'b00100101;
			21: led = 8'b10011111;
			21: led2 = 8'b00100101;
			22: led = 8'b00100101;
			22: led2 = 8'b00100101;
			23: led = 8'b00001101;
			23: led2 = 8'b00100101;
			24: led = 8'b10011001;
			24: led2 = 8'b00100101;
			25: led = 8'b01001001;
			25: led2 = 8'b00100101;
			26: led = 8'b01000001;
			26: led2 = 8'b00100101;
			27: led = 8'b00011111;
			27: led2 = 8'b00100101;
			28: led = 8'b00000001;
			28: led2 = 8'b00100101;
			29: led = 8'b00001001;
			29: led2 = 8'b00100101;
			
			
			30: led = 8'b00000011;
	   	30: led2 = 8'b00001101;
			31: led = 8'b10011111;
			31: led2 = 8'b00001101;
			32: led = 8'b00100101;
			32: led2 = 8'b00001101;
			33: led = 8'b00001101;
			33: led2 = 8'b00001101;
			34: led = 8'b10011001;
			34: led2 = 8'b00001101;
			35: led = 8'b01001001;
			35: led2 = 8'b00001101;
			36: led = 8'b01000001;
			36: led2 = 8'b00001101;
			37: led = 8'b00011111;
			37: led2 = 8'b00001101;
			38: led = 8'b00000001;
			38: led2 = 8'b00001101;
			39: led = 8'b00001001;
			39: led2 = 8'b00001101;
			
			default: led = 8'b11111111;
			
		endcase
		

endmodule
